`define KNN_ADDR_W 3  //address width
`define KNN_WDATA_W 128 //write data width (32 * 4)
`ifndef DATA_W
 `define DATA_W 32      //cpu data width
`endif
